
--------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_wait_pkg_v1 IS

COMPONENT ccs_in_wait_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    rdy    : OUT std_logic;
    ivld   : OUT std_logic;
    dat    : IN  std_logic_vector(width-1 DOWNTO 0);
    irdy   : IN  std_logic;
    vld    : IN  std_logic
   );
END COMPONENT;

END ccs_in_wait_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_wait_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    rdy   : OUT std_logic;
    ivld  : OUT std_logic;
    dat   : IN  std_logic_vector(width-1 DOWNTO 0);
    irdy  : IN  std_logic;
    vld   : IN  std_logic
  );
END ccs_in_wait_v1;

ARCHITECTURE beh OF ccs_in_wait_v1 IS
  constant stall_const : std_logic := '0';
  SIGNAL stall_ctrl : std_logic;
BEGIN
  stall_ctrl <= stall_const;

  idat <= dat;
  rdy  <= irdy and not stall_ctrl;
  ivld <= vld and not stall_ctrl;

END beh;


--------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_out_wait_pkg_v1 IS

COMPONENT ccs_out_wait_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    dat    : OUT std_logic_vector(width-1 DOWNTO 0);
    irdy   : OUT std_logic;
    vld    : OUT std_logic;
    idat   : IN  std_logic_vector(width-1 DOWNTO 0);
    rdy    : IN  std_logic;
    ivld   : IN  std_logic
  );
END COMPONENT;

END ccs_out_wait_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_out_wait_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    dat   : OUT std_logic_vector(width-1 DOWNTO 0);
    irdy  : OUT std_logic;
    vld   : OUT std_logic;
    idat  : IN  std_logic_vector(width-1 DOWNTO 0);
    rdy   : IN  std_logic;
    ivld  : IN  std_logic
  );
END ccs_out_wait_v1;

ARCHITECTURE beh OF ccs_out_wait_v1 IS
  constant stall_const : std_logic := '0';
  SIGNAL stall_ctrl : std_logic;
BEGIN
  stall_ctrl <= stall_const;

  dat  <= idat;
  irdy <= rdy and not stall_ctrl;
  vld  <= ivld and not stall_ctrl;

END beh;


--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2023.2/1059873 Production Release
--  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
-- 
--  Generated by:   r12016@cad40
--  Generated date: Sun Mar 24 17:31:51 2024
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    fir_run_run_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_run_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    run_wen : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END fir_run_run_fsm;

ARCHITECTURE v2 OF fir_run_run_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for fir_run_run_fsm_1
  TYPE fir_run_run_fsm_1_ST IS (run_rlp_C_0, main_C_0);

  SIGNAL state_var : fir_run_run_fsm_1_ST;
  SIGNAL state_var_NS : fir_run_run_fsm_1_ST;

BEGIN
  fir_run_run_fsm_1 : PROCESS (state_var)
  BEGIN
    CASE state_var IS
      WHEN main_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10");
        state_var_NS <= main_C_0;
      -- run_rlp_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "01");
        state_var_NS <= main_C_0;
    END CASE;
  END PROCESS fir_run_run_fsm_1;

  fir_run_run_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= run_rlp_C_0;
      ELSE
        IF ( run_wen = '1' ) THEN
          state_var <= state_var_NS;
        END IF;
      END IF;
    END IF;
  END PROCESS fir_run_run_fsm_1_REG;

END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run_staller
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_staller IS
  PORT(
    run_wen : OUT STD_LOGIC;
    input_rsci_wen_comp : IN STD_LOGIC;
    output_rsci_wen_comp : IN STD_LOGIC
  );
END fir_run_staller;

ARCHITECTURE v2 OF fir_run_staller IS
  -- Default Constants

BEGIN
  run_wen <= input_rsci_wen_comp AND output_rsci_wen_comp;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run_output_rsci_output_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_output_rsci_output_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    output_rsci_oswt : IN STD_LOGIC;
    output_rsci_wen_comp : OUT STD_LOGIC;
    output_rsci_biwt : IN STD_LOGIC;
    output_rsci_bdwt : IN STD_LOGIC;
    output_rsci_bcwt : OUT STD_LOGIC
  );
END fir_run_output_rsci_output_wait_dp;

ARCHITECTURE v2 OF fir_run_output_rsci_output_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL output_rsci_bcwt_drv : STD_LOGIC;

BEGIN
  -- Output Reader Assignments
  output_rsci_bcwt <= output_rsci_bcwt_drv;

  output_rsci_wen_comp <= (NOT output_rsci_oswt) OR output_rsci_biwt OR output_rsci_bcwt_drv;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_bcwt_drv <= '0';
      ELSE
        output_rsci_bcwt_drv <= NOT((NOT(output_rsci_bcwt_drv OR output_rsci_biwt))
            OR output_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run_output_rsci_output_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_output_rsci_output_wait_ctrl IS
  PORT(
    run_wen : IN STD_LOGIC;
    output_rsci_oswt : IN STD_LOGIC;
    output_rsci_biwt : OUT STD_LOGIC;
    output_rsci_bdwt : OUT STD_LOGIC;
    output_rsci_bcwt : IN STD_LOGIC;
    output_rsci_irdy : IN STD_LOGIC;
    output_rsci_ivld_run_sct : OUT STD_LOGIC
  );
END fir_run_output_rsci_output_wait_ctrl;

ARCHITECTURE v2 OF fir_run_output_rsci_output_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL output_rsci_ogwt : STD_LOGIC;

BEGIN
  output_rsci_bdwt <= output_rsci_oswt AND run_wen;
  output_rsci_biwt <= output_rsci_ogwt AND output_rsci_irdy;
  output_rsci_ogwt <= output_rsci_oswt AND (NOT output_rsci_bcwt);
  output_rsci_ivld_run_sct <= output_rsci_ogwt;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run_input_rsci_input_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_input_rsci_input_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsci_oswt : IN STD_LOGIC;
    input_rsci_wen_comp : OUT STD_LOGIC;
    input_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    input_rsci_biwt : IN STD_LOGIC;
    input_rsci_bdwt : IN STD_LOGIC;
    input_rsci_bcwt : OUT STD_LOGIC;
    input_rsci_idat : IN STD_LOGIC_VECTOR (7 DOWNTO 0)
  );
END fir_run_input_rsci_input_wait_dp;

ARCHITECTURE v2 OF fir_run_input_rsci_input_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL input_rsci_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL input_rsci_idat_bfwt : STD_LOGIC_VECTOR (7 DOWNTO 0);

  FUNCTION MUX_v_8_2_2(input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  input_rsci_bcwt <= input_rsci_bcwt_drv;

  input_rsci_wen_comp <= (NOT input_rsci_oswt) OR input_rsci_biwt OR input_rsci_bcwt_drv;
  input_rsci_idat_mxwt <= MUX_v_8_2_2(input_rsci_idat, input_rsci_idat_bfwt, input_rsci_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        input_rsci_bcwt_drv <= '0';
      ELSE
        input_rsci_bcwt_drv <= NOT((NOT(input_rsci_bcwt_drv OR input_rsci_biwt))
            OR input_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        input_rsci_idat_bfwt <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( input_rsci_biwt = '1' ) THEN
        input_rsci_idat_bfwt <= input_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run_input_rsci_input_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_input_rsci_input_wait_ctrl IS
  PORT(
    run_wen : IN STD_LOGIC;
    input_rsci_oswt : IN STD_LOGIC;
    input_rsci_biwt : OUT STD_LOGIC;
    input_rsci_bdwt : OUT STD_LOGIC;
    input_rsci_bcwt : IN STD_LOGIC;
    input_rsci_irdy_run_sct : OUT STD_LOGIC;
    input_rsci_ivld : IN STD_LOGIC
  );
END fir_run_input_rsci_input_wait_ctrl;

ARCHITECTURE v2 OF fir_run_input_rsci_input_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL input_rsci_ogwt : STD_LOGIC;

BEGIN
  input_rsci_bdwt <= input_rsci_oswt AND run_wen;
  input_rsci_biwt <= input_rsci_ogwt AND input_rsci_ivld;
  input_rsci_ogwt <= input_rsci_oswt AND (NOT input_rsci_bcwt);
  input_rsci_irdy_run_sct <= input_rsci_ogwt;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator_run_run_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator_run_run_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    run_wen : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
  );
END decimator_run_run_fsm;

ARCHITECTURE v2 OF decimator_run_run_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for decimator_run_run_fsm_1
  TYPE decimator_run_run_fsm_1_ST IS (run_rlp_C_0, main_C_0, main_C_1);

  SIGNAL state_var : decimator_run_run_fsm_1_ST;
  SIGNAL state_var_NS : decimator_run_run_fsm_1_ST;

BEGIN
  decimator_run_run_fsm_1 : PROCESS (state_var)
  BEGIN
    CASE state_var IS
      WHEN main_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010");
        state_var_NS <= main_C_1;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100");
        state_var_NS <= main_C_0;
      -- run_rlp_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "001");
        state_var_NS <= main_C_0;
    END CASE;
  END PROCESS decimator_run_run_fsm_1;

  decimator_run_run_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= run_rlp_C_0;
      ELSE
        IF ( run_wen = '1' ) THEN
          state_var <= state_var_NS;
        END IF;
      END IF;
    END IF;
  END PROCESS decimator_run_run_fsm_1_REG;

END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator_run_staller
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator_run_staller IS
  PORT(
    run_wen : OUT STD_LOGIC;
    din_rsci_wen_comp : IN STD_LOGIC;
    dout_rsci_wen_comp : IN STD_LOGIC
  );
END decimator_run_staller;

ARCHITECTURE v2 OF decimator_run_staller IS
  -- Default Constants

BEGIN
  run_wen <= din_rsci_wen_comp AND dout_rsci_wen_comp;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator_run_dout_rsci_dout_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator_run_dout_rsci_dout_wait_ctrl IS
  PORT(
    dout_rsci_iswt0 : IN STD_LOGIC;
    dout_rsci_biwt : OUT STD_LOGIC;
    dout_rsci_irdy : IN STD_LOGIC
  );
END decimator_run_dout_rsci_dout_wait_ctrl;

ARCHITECTURE v2 OF decimator_run_dout_rsci_dout_wait_ctrl IS
  -- Default Constants

BEGIN
  dout_rsci_biwt <= dout_rsci_iswt0 AND dout_rsci_irdy;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator_run_din_rsci_din_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator_run_din_rsci_din_wait_ctrl IS
  PORT(
    din_rsci_iswt0 : IN STD_LOGIC;
    din_rsci_biwt : OUT STD_LOGIC;
    din_rsci_ivld : IN STD_LOGIC
  );
END decimator_run_din_rsci_din_wait_ctrl;

ARCHITECTURE v2 OF decimator_run_din_rsci_din_wait_ctrl IS
  -- Default Constants

BEGIN
  din_rsci_biwt <= din_rsci_iswt0 AND din_rsci_ivld;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run_output_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_output_rsci IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    output_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    output_rsc_vld : OUT STD_LOGIC;
    output_rsc_rdy : IN STD_LOGIC;
    run_wen : IN STD_LOGIC;
    output_rsci_oswt : IN STD_LOGIC;
    output_rsci_wen_comp : OUT STD_LOGIC;
    output_rsci_idat : IN STD_LOGIC_VECTOR (7 DOWNTO 0)
  );
END fir_run_output_rsci;

ARCHITECTURE v2 OF fir_run_output_rsci IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL output_rsci_biwt : STD_LOGIC;
  SIGNAL output_rsci_bdwt : STD_LOGIC;
  SIGNAL output_rsci_bcwt : STD_LOGIC;
  SIGNAL output_rsci_irdy : STD_LOGIC;
  SIGNAL output_rsci_ivld_run_sct : STD_LOGIC;

  SIGNAL output_rsci_idat_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL output_rsci_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);

  COMPONENT fir_run_output_rsci_output_wait_ctrl
    PORT(
      run_wen : IN STD_LOGIC;
      output_rsci_oswt : IN STD_LOGIC;
      output_rsci_biwt : OUT STD_LOGIC;
      output_rsci_bdwt : OUT STD_LOGIC;
      output_rsci_bcwt : IN STD_LOGIC;
      output_rsci_irdy : IN STD_LOGIC;
      output_rsci_ivld_run_sct : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT fir_run_output_rsci_output_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      output_rsci_oswt : IN STD_LOGIC;
      output_rsci_wen_comp : OUT STD_LOGIC;
      output_rsci_biwt : IN STD_LOGIC;
      output_rsci_bdwt : IN STD_LOGIC;
      output_rsci_bcwt : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  output_rsci : work.ccs_out_wait_pkg_v1.ccs_out_wait_v1
    GENERIC MAP(
      rscid => 3,
      width => 8
      )
    PORT MAP(
      irdy => output_rsci_irdy,
      ivld => output_rsci_ivld_run_sct,
      idat => output_rsci_idat_1,
      rdy => output_rsc_rdy,
      vld => output_rsc_vld,
      dat => output_rsci_dat
    );
  output_rsci_idat_1 <= output_rsci_idat;
  output_rsc_dat <= output_rsci_dat;

  fir_run_output_rsci_output_wait_ctrl_inst : fir_run_output_rsci_output_wait_ctrl
    PORT MAP(
      run_wen => run_wen,
      output_rsci_oswt => output_rsci_oswt,
      output_rsci_biwt => output_rsci_biwt,
      output_rsci_bdwt => output_rsci_bdwt,
      output_rsci_bcwt => output_rsci_bcwt,
      output_rsci_irdy => output_rsci_irdy,
      output_rsci_ivld_run_sct => output_rsci_ivld_run_sct
    );
  fir_run_output_rsci_output_wait_dp_inst : fir_run_output_rsci_output_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      output_rsci_oswt => output_rsci_oswt,
      output_rsci_wen_comp => output_rsci_wen_comp,
      output_rsci_biwt => output_rsci_biwt,
      output_rsci_bdwt => output_rsci_bdwt,
      output_rsci_bcwt => output_rsci_bcwt
    );
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run_input_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run_input_rsci IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    input_rsc_vld : IN STD_LOGIC;
    input_rsc_rdy : OUT STD_LOGIC;
    run_wen : IN STD_LOGIC;
    input_rsci_oswt : IN STD_LOGIC;
    input_rsci_wen_comp : OUT STD_LOGIC;
    input_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
  );
END fir_run_input_rsci;

ARCHITECTURE v2 OF fir_run_input_rsci IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL input_rsci_biwt : STD_LOGIC;
  SIGNAL input_rsci_bdwt : STD_LOGIC;
  SIGNAL input_rsci_bcwt : STD_LOGIC;
  SIGNAL input_rsci_irdy_run_sct : STD_LOGIC;
  SIGNAL input_rsci_ivld : STD_LOGIC;
  SIGNAL input_rsci_idat : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL input_rsci_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL input_rsci_idat_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);

  COMPONENT fir_run_input_rsci_input_wait_ctrl
    PORT(
      run_wen : IN STD_LOGIC;
      input_rsci_oswt : IN STD_LOGIC;
      input_rsci_biwt : OUT STD_LOGIC;
      input_rsci_bdwt : OUT STD_LOGIC;
      input_rsci_bcwt : IN STD_LOGIC;
      input_rsci_irdy_run_sct : OUT STD_LOGIC;
      input_rsci_ivld : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT fir_run_input_rsci_input_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      input_rsci_oswt : IN STD_LOGIC;
      input_rsci_wen_comp : OUT STD_LOGIC;
      input_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      input_rsci_biwt : IN STD_LOGIC;
      input_rsci_bdwt : IN STD_LOGIC;
      input_rsci_bcwt : OUT STD_LOGIC;
      input_rsci_idat : IN STD_LOGIC_VECTOR (7 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL fir_run_input_rsci_input_wait_dp_inst_input_rsci_idat_mxwt : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL fir_run_input_rsci_input_wait_dp_inst_input_rsci_idat : STD_LOGIC_VECTOR
      (7 DOWNTO 0);

BEGIN
  input_rsci : work.ccs_in_wait_pkg_v1.ccs_in_wait_v1
    GENERIC MAP(
      rscid => 1,
      width => 8
      )
    PORT MAP(
      rdy => input_rsc_rdy,
      vld => input_rsc_vld,
      dat => input_rsci_dat,
      irdy => input_rsci_irdy_run_sct,
      ivld => input_rsci_ivld,
      idat => input_rsci_idat_1
    );
  input_rsci_dat <= input_rsc_dat;
  input_rsci_idat <= input_rsci_idat_1;

  fir_run_input_rsci_input_wait_ctrl_inst : fir_run_input_rsci_input_wait_ctrl
    PORT MAP(
      run_wen => run_wen,
      input_rsci_oswt => input_rsci_oswt,
      input_rsci_biwt => input_rsci_biwt,
      input_rsci_bdwt => input_rsci_bdwt,
      input_rsci_bcwt => input_rsci_bcwt,
      input_rsci_irdy_run_sct => input_rsci_irdy_run_sct,
      input_rsci_ivld => input_rsci_ivld
    );
  fir_run_input_rsci_input_wait_dp_inst : fir_run_input_rsci_input_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      input_rsci_oswt => input_rsci_oswt,
      input_rsci_wen_comp => input_rsci_wen_comp,
      input_rsci_idat_mxwt => fir_run_input_rsci_input_wait_dp_inst_input_rsci_idat_mxwt,
      input_rsci_biwt => input_rsci_biwt,
      input_rsci_bdwt => input_rsci_bdwt,
      input_rsci_bcwt => input_rsci_bcwt,
      input_rsci_idat => fir_run_input_rsci_input_wait_dp_inst_input_rsci_idat
    );
  input_rsci_idat_mxwt <= fir_run_input_rsci_input_wait_dp_inst_input_rsci_idat_mxwt;
  fir_run_input_rsci_input_wait_dp_inst_input_rsci_idat <= input_rsci_idat;

END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator_run_dout_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator_run_dout_rsci IS
  PORT(
    dout_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    dout_rsc_vld : OUT STD_LOGIC;
    dout_rsc_rdy : IN STD_LOGIC;
    dout_rsci_oswt : IN STD_LOGIC;
    dout_rsci_wen_comp : OUT STD_LOGIC;
    dout_rsci_idat : IN STD_LOGIC_VECTOR (7 DOWNTO 0)
  );
END decimator_run_dout_rsci;

ARCHITECTURE v2 OF decimator_run_dout_rsci IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL dout_rsci_biwt : STD_LOGIC;
  SIGNAL dout_rsci_irdy : STD_LOGIC;

  SIGNAL dout_rsci_idat_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL dout_rsci_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);

  COMPONENT decimator_run_dout_rsci_dout_wait_ctrl
    PORT(
      dout_rsci_iswt0 : IN STD_LOGIC;
      dout_rsci_biwt : OUT STD_LOGIC;
      dout_rsci_irdy : IN STD_LOGIC
    );
  END COMPONENT;
BEGIN
  dout_rsci : work.ccs_out_wait_pkg_v1.ccs_out_wait_v1
    GENERIC MAP(
      rscid => 6,
      width => 8
      )
    PORT MAP(
      irdy => dout_rsci_irdy,
      ivld => dout_rsci_oswt,
      idat => dout_rsci_idat_1,
      rdy => dout_rsc_rdy,
      vld => dout_rsc_vld,
      dat => dout_rsci_dat
    );
  dout_rsci_idat_1 <= dout_rsci_idat;
  dout_rsc_dat <= dout_rsci_dat;

  decimator_run_dout_rsci_dout_wait_ctrl_inst : decimator_run_dout_rsci_dout_wait_ctrl
    PORT MAP(
      dout_rsci_iswt0 => dout_rsci_oswt,
      dout_rsci_biwt => dout_rsci_biwt,
      dout_rsci_irdy => dout_rsci_irdy
    );
  dout_rsci_wen_comp <= (NOT dout_rsci_oswt) OR dout_rsci_biwt;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator_run_din_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator_run_din_rsci IS
  PORT(
    din_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    din_rsc_vld : IN STD_LOGIC;
    din_rsc_rdy : OUT STD_LOGIC;
    din_rsci_oswt : IN STD_LOGIC;
    din_rsci_wen_comp : OUT STD_LOGIC;
    din_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
  );
END decimator_run_din_rsci;

ARCHITECTURE v2 OF decimator_run_din_rsci IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL din_rsci_biwt : STD_LOGIC;
  SIGNAL din_rsci_ivld : STD_LOGIC;
  SIGNAL din_rsci_idat : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL din_rsci_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL din_rsci_idat_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);

  COMPONENT decimator_run_din_rsci_din_wait_ctrl
    PORT(
      din_rsci_iswt0 : IN STD_LOGIC;
      din_rsci_biwt : OUT STD_LOGIC;
      din_rsci_ivld : IN STD_LOGIC
    );
  END COMPONENT;
BEGIN
  din_rsci : work.ccs_in_wait_pkg_v1.ccs_in_wait_v1
    GENERIC MAP(
      rscid => 5,
      width => 8
      )
    PORT MAP(
      rdy => din_rsc_rdy,
      vld => din_rsc_vld,
      dat => din_rsci_dat,
      irdy => din_rsci_oswt,
      ivld => din_rsci_ivld,
      idat => din_rsci_idat_1
    );
  din_rsci_dat <= din_rsc_dat;
  din_rsci_idat <= din_rsci_idat_1;

  decimator_run_din_rsci_din_wait_ctrl_inst : decimator_run_din_rsci_din_wait_ctrl
    PORT MAP(
      din_rsci_iswt0 => din_rsci_oswt,
      din_rsci_biwt => din_rsci_biwt,
      din_rsci_ivld => din_rsci_ivld
    );
  din_rsci_idat_mxwt <= din_rsci_idat;
  din_rsci_wen_comp <= (NOT din_rsci_oswt) OR din_rsci_biwt;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir_run
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir_run IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    input_rsc_vld : IN STD_LOGIC;
    input_rsc_rdy : OUT STD_LOGIC;
    coeffs : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    output_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    output_rsc_vld : OUT STD_LOGIC;
    output_rsc_rdy : IN STD_LOGIC
  );
END fir_run;

ARCHITECTURE v2 OF fir_run IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL run_wen : STD_LOGIC;
  SIGNAL input_rsci_wen_comp : STD_LOGIC;
  SIGNAL input_rsci_idat_mxwt : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL output_rsci_wen_comp : STD_LOGIC;
  SIGNAL output_rsci_idat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reg_output_rsci_iswt0_cse : STD_LOGIC;
  SIGNAL reg_input_rsci_iswt0_cse : STD_LOGIC;
  SIGNAL and_18_cse : STD_LOGIC;
  SIGNAL regs_1_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL regs_0_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL MAC_asn_4_itm : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL MAC_asn_8_itm : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL MAC_asn_10_itm : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL MAC_asn_12_itm : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL MAC_asn_14_itm : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL MAC_8_acc_1_nl : STD_LOGIC_VECTOR (18 DOWNTO 0);
  SIGNAL MAC_3_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_4_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_7_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_8_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_5_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_6_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_1_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_2_mul_nl : STD_LOGIC_VECTOR (15 DOWNTO 0);
  COMPONENT fir_run_input_rsci
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      input_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      input_rsc_vld : IN STD_LOGIC;
      input_rsc_rdy : OUT STD_LOGIC;
      run_wen : IN STD_LOGIC;
      input_rsci_oswt : IN STD_LOGIC;
      input_rsci_wen_comp : OUT STD_LOGIC;
      input_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL fir_run_input_rsci_inst_input_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL fir_run_input_rsci_inst_input_rsci_idat_mxwt : STD_LOGIC_VECTOR (7 DOWNTO
      0);

  COMPONENT fir_run_output_rsci
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      output_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      output_rsc_vld : OUT STD_LOGIC;
      output_rsc_rdy : IN STD_LOGIC;
      run_wen : IN STD_LOGIC;
      output_rsci_oswt : IN STD_LOGIC;
      output_rsci_wen_comp : OUT STD_LOGIC;
      output_rsci_idat : IN STD_LOGIC_VECTOR (7 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL fir_run_output_rsci_inst_output_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL fir_run_output_rsci_inst_output_rsci_idat : STD_LOGIC_VECTOR (7 DOWNTO 0);

  COMPONENT fir_run_staller
    PORT(
      run_wen : OUT STD_LOGIC;
      input_rsci_wen_comp : IN STD_LOGIC;
      output_rsci_wen_comp : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT fir_run_run_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      run_wen : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL fir_run_run_fsm_inst_fsm_output : STD_LOGIC_VECTOR (1 DOWNTO 0);

BEGIN
  fir_run_input_rsci_inst : fir_run_input_rsci
    PORT MAP(
      clk => clk,
      rst => rst,
      input_rsc_dat => fir_run_input_rsci_inst_input_rsc_dat,
      input_rsc_vld => input_rsc_vld,
      input_rsc_rdy => input_rsc_rdy,
      run_wen => run_wen,
      input_rsci_oswt => reg_input_rsci_iswt0_cse,
      input_rsci_wen_comp => input_rsci_wen_comp,
      input_rsci_idat_mxwt => fir_run_input_rsci_inst_input_rsci_idat_mxwt
    );
  fir_run_input_rsci_inst_input_rsc_dat <= input_rsc_dat;
  input_rsci_idat_mxwt <= fir_run_input_rsci_inst_input_rsci_idat_mxwt;

  fir_run_output_rsci_inst : fir_run_output_rsci
    PORT MAP(
      clk => clk,
      rst => rst,
      output_rsc_dat => fir_run_output_rsci_inst_output_rsc_dat,
      output_rsc_vld => output_rsc_vld,
      output_rsc_rdy => output_rsc_rdy,
      run_wen => run_wen,
      output_rsci_oswt => reg_output_rsci_iswt0_cse,
      output_rsci_wen_comp => output_rsci_wen_comp,
      output_rsci_idat => fir_run_output_rsci_inst_output_rsci_idat
    );
  output_rsc_dat <= fir_run_output_rsci_inst_output_rsc_dat;
  fir_run_output_rsci_inst_output_rsci_idat <= output_rsci_idat;

  fir_run_staller_inst : fir_run_staller
    PORT MAP(
      run_wen => run_wen,
      input_rsci_wen_comp => input_rsci_wen_comp,
      output_rsci_wen_comp => output_rsci_wen_comp
    );
  fir_run_run_fsm_inst : fir_run_run_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      run_wen => run_wen,
      fsm_output => fir_run_run_fsm_inst_fsm_output
    );
  fsm_output <= fir_run_run_fsm_inst_fsm_output;

  and_18_cse <= run_wen AND (NOT (fsm_output(0)));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        output_rsci_idat <= STD_LOGIC_VECTOR'( "00000000");
        regs_0_sva <= STD_LOGIC_VECTOR'( "00000000");
        MAC_asn_4_itm <= STD_LOGIC_VECTOR'( "00000000");
        regs_1_sva <= STD_LOGIC_VECTOR'( "00000000");
        MAC_asn_8_itm <= STD_LOGIC_VECTOR'( "00000000");
        MAC_asn_10_itm <= STD_LOGIC_VECTOR'( "00000000");
        MAC_asn_12_itm <= STD_LOGIC_VECTOR'( "00000000");
        MAC_asn_14_itm <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( and_18_cse = '1' ) THEN
        output_rsci_idat <= MAC_8_acc_1_nl(18 DOWNTO 11);
        regs_0_sva <= input_rsci_idat_mxwt;
        MAC_asn_4_itm <= regs_1_sva;
        regs_1_sva <= regs_0_sva;
        MAC_asn_8_itm <= MAC_asn_10_itm;
        MAC_asn_10_itm <= MAC_asn_4_itm;
        MAC_asn_12_itm <= MAC_asn_14_itm;
        MAC_asn_14_itm <= MAC_asn_8_itm;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_output_rsci_iswt0_cse <= '0';
        reg_input_rsci_iswt0_cse <= '0';
      ELSIF ( run_wen = '1' ) THEN
        reg_output_rsci_iswt0_cse <= fsm_output(1);
        reg_input_rsci_iswt0_cse <= '1';
      END IF;
    END IF;
  END PROCESS;
  MAC_3_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(47 DOWNTO 40))
      * SIGNED(MAC_asn_8_itm)), 16));
  MAC_4_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(39 DOWNTO 32))
      * SIGNED(MAC_asn_10_itm)), 16));
  MAC_7_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(15 DOWNTO 8))
      * SIGNED(regs_0_sva)), 16));
  MAC_8_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(7 DOWNTO 0))
      * SIGNED(input_rsci_idat_mxwt)), 16));
  MAC_5_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(31 DOWNTO 24))
      * SIGNED(MAC_asn_4_itm)), 16));
  MAC_6_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(23 DOWNTO 16))
      * SIGNED(regs_1_sva)), 16));
  MAC_1_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(63 DOWNTO 56))
      * SIGNED(MAC_asn_12_itm)), 16));
  MAC_2_mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(coeffs(55 DOWNTO 48))
      * SIGNED(MAC_asn_14_itm)), 16));
  MAC_8_acc_1_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(SIGNED(MAC_3_mul_nl),
      19) + CONV_SIGNED(SIGNED(MAC_4_mul_nl), 19) + CONV_SIGNED(SIGNED(MAC_7_mul_nl),
      19) + CONV_SIGNED(SIGNED(MAC_8_mul_nl), 19) + CONV_SIGNED(SIGNED(MAC_5_mul_nl),
      19) + CONV_SIGNED(SIGNED(MAC_6_mul_nl), 19) + CONV_SIGNED(SIGNED(MAC_1_mul_nl),
      19) + CONV_SIGNED(SIGNED(MAC_2_mul_nl), 19), 19));
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator_run
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator_run IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    din_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    din_rsc_vld : IN STD_LOGIC;
    din_rsc_rdy : OUT STD_LOGIC;
    dout_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    dout_rsc_vld : OUT STD_LOGIC;
    dout_rsc_rdy : IN STD_LOGIC
  );
END decimator_run;

ARCHITECTURE v2 OF decimator_run IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL run_wen : STD_LOGIC;
  SIGNAL din_rsci_wen_comp : STD_LOGIC;
  SIGNAL din_rsci_idat_mxwt : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL dout_rsci_wen_comp : STD_LOGIC;
  SIGNAL dout_rsci_idat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL equal_tmp : STD_LOGIC;
  SIGNAL reg_dout_rsci_iswt0_cse : STD_LOGIC;
  SIGNAL reg_din_rsci_iswt0_cse : STD_LOGIC;
  SIGNAL count_2_0_sva_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT decimator_run_din_rsci
    PORT(
      din_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      din_rsc_vld : IN STD_LOGIC;
      din_rsc_rdy : OUT STD_LOGIC;
      din_rsci_oswt : IN STD_LOGIC;
      din_rsci_wen_comp : OUT STD_LOGIC;
      din_rsci_idat_mxwt : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL decimator_run_din_rsci_inst_din_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL decimator_run_din_rsci_inst_din_rsci_idat_mxwt : STD_LOGIC_VECTOR (7 DOWNTO
      0);

  COMPONENT decimator_run_dout_rsci
    PORT(
      dout_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      dout_rsc_vld : OUT STD_LOGIC;
      dout_rsc_rdy : IN STD_LOGIC;
      dout_rsci_oswt : IN STD_LOGIC;
      dout_rsci_wen_comp : OUT STD_LOGIC;
      dout_rsci_idat : IN STD_LOGIC_VECTOR (7 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL decimator_run_dout_rsci_inst_dout_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL decimator_run_dout_rsci_inst_dout_rsci_idat : STD_LOGIC_VECTOR (7 DOWNTO
      0);

  COMPONENT decimator_run_staller
    PORT(
      run_wen : OUT STD_LOGIC;
      din_rsci_wen_comp : IN STD_LOGIC;
      dout_rsci_wen_comp : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT decimator_run_run_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      run_wen : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL decimator_run_run_fsm_inst_fsm_output : STD_LOGIC_VECTOR (2 DOWNTO 0);

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

BEGIN
  decimator_run_din_rsci_inst : decimator_run_din_rsci
    PORT MAP(
      din_rsc_dat => decimator_run_din_rsci_inst_din_rsc_dat,
      din_rsc_vld => din_rsc_vld,
      din_rsc_rdy => din_rsc_rdy,
      din_rsci_oswt => reg_din_rsci_iswt0_cse,
      din_rsci_wen_comp => din_rsci_wen_comp,
      din_rsci_idat_mxwt => decimator_run_din_rsci_inst_din_rsci_idat_mxwt
    );
  decimator_run_din_rsci_inst_din_rsc_dat <= din_rsc_dat;
  din_rsci_idat_mxwt <= decimator_run_din_rsci_inst_din_rsci_idat_mxwt;

  decimator_run_dout_rsci_inst : decimator_run_dout_rsci
    PORT MAP(
      dout_rsc_dat => decimator_run_dout_rsci_inst_dout_rsc_dat,
      dout_rsc_vld => dout_rsc_vld,
      dout_rsc_rdy => dout_rsc_rdy,
      dout_rsci_oswt => reg_dout_rsci_iswt0_cse,
      dout_rsci_wen_comp => dout_rsci_wen_comp,
      dout_rsci_idat => decimator_run_dout_rsci_inst_dout_rsci_idat
    );
  dout_rsc_dat <= decimator_run_dout_rsci_inst_dout_rsc_dat;
  decimator_run_dout_rsci_inst_dout_rsci_idat <= dout_rsci_idat;

  decimator_run_staller_inst : decimator_run_staller
    PORT MAP(
      run_wen => run_wen,
      din_rsci_wen_comp => din_rsci_wen_comp,
      dout_rsci_wen_comp => dout_rsci_wen_comp
    );
  decimator_run_run_fsm_inst : decimator_run_run_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      run_wen => run_wen,
      fsm_output => decimator_run_run_fsm_inst_fsm_output
    );
  fsm_output <= decimator_run_run_fsm_inst_fsm_output;

  equal_tmp <= NOT(CONV_SL_1_1(count_2_0_sva_1_0/=STD_LOGIC_VECTOR'("00")));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        dout_rsci_idat <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (run_wen AND equal_tmp AND (fsm_output(1))) = '1' ) THEN
        dout_rsci_idat <= din_rsci_idat_mxwt;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_dout_rsci_iswt0_cse <= '0';
        reg_din_rsci_iswt0_cse <= '0';
      ELSIF ( run_wen = '1' ) THEN
        reg_dout_rsci_iswt0_cse <= equal_tmp AND (fsm_output(1));
        reg_din_rsci_iswt0_cse <= NOT (fsm_output(1));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        count_2_0_sva_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (run_wen AND (fsm_output(1))) = '1' ) THEN
        count_2_0_sva_1_0 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(count_2_0_sva_1_0)
            + SIGNED'( "01"), 2));
      END IF;
    END IF;
  END PROCESS;
END v2;

-- ------------------------------------------------------------------
--  Design Unit:    fir
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY fir IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    input_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    input_rsc_vld : IN STD_LOGIC;
    input_rsc_rdy : OUT STD_LOGIC;
    coeffs : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    output_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    output_rsc_vld : OUT STD_LOGIC;
    output_rsc_rdy : IN STD_LOGIC
  );
END fir;

ARCHITECTURE v2 OF fir IS
  -- Default Constants

  COMPONENT fir_run
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      input_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      input_rsc_vld : IN STD_LOGIC;
      input_rsc_rdy : OUT STD_LOGIC;
      coeffs : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      output_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      output_rsc_vld : OUT STD_LOGIC;
      output_rsc_rdy : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL fir_run_inst_input_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL fir_run_inst_coeffs : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL fir_run_inst_output_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);

BEGIN
  fir_run_inst : fir_run
    PORT MAP(
      clk => clk,
      rst => rst,
      input_rsc_dat => fir_run_inst_input_rsc_dat,
      input_rsc_vld => input_rsc_vld,
      input_rsc_rdy => input_rsc_rdy,
      coeffs => fir_run_inst_coeffs,
      output_rsc_dat => fir_run_inst_output_rsc_dat,
      output_rsc_vld => output_rsc_vld,
      output_rsc_rdy => output_rsc_rdy
    );
  fir_run_inst_input_rsc_dat <= input_rsc_dat;
  fir_run_inst_coeffs <= coeffs;
  output_rsc_dat <= fir_run_inst_output_rsc_dat;

END v2;

-- ------------------------------------------------------------------
--  Design Unit:    decimator
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY decimator IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    din_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    din_rsc_vld : IN STD_LOGIC;
    din_rsc_rdy : OUT STD_LOGIC;
    dout_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    dout_rsc_vld : OUT STD_LOGIC;
    dout_rsc_rdy : IN STD_LOGIC
  );
END decimator;

ARCHITECTURE v2 OF decimator IS
  -- Default Constants

  COMPONENT decimator_run
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      din_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      din_rsc_vld : IN STD_LOGIC;
      din_rsc_rdy : OUT STD_LOGIC;
      dout_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      dout_rsc_vld : OUT STD_LOGIC;
      dout_rsc_rdy : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL decimator_run_inst_din_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL decimator_run_inst_dout_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);

BEGIN
  decimator_run_inst : decimator_run
    PORT MAP(
      clk => clk,
      rst => rst,
      din_rsc_dat => decimator_run_inst_din_rsc_dat,
      din_rsc_vld => din_rsc_vld,
      din_rsc_rdy => din_rsc_rdy,
      dout_rsc_dat => decimator_run_inst_dout_rsc_dat,
      dout_rsc_vld => dout_rsc_vld,
      dout_rsc_rdy => dout_rsc_rdy
    );
  decimator_run_inst_din_rsc_dat <= din_rsc_dat;
  dout_rsc_dat <= decimator_run_inst_dout_rsc_dat;

END v2;

-- ------------------------------------------------------------------
--  Design Unit:    top
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_wait_pkg_v1.ALL;
USE work.ccs_out_wait_pkg_v1.ALL;


ENTITY top IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    din_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    din_rsc_vld : IN STD_LOGIC;
    din_rsc_rdy : OUT STD_LOGIC;
    coeffs : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    dout_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    dout_rsc_vld : OUT STD_LOGIC;
    dout_rsc_rdy : IN STD_LOGIC
  );
END top;

ARCHITECTURE v2 OF top IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL output_rsc_dat_n_block0 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL output_rsc_dat_n_block1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL dout_rsc_dat_n_block2 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL input_rsc_rdy_n_block0_bud : STD_LOGIC;
  SIGNAL output_rsc_vld_n_block0_bud : STD_LOGIC;
  SIGNAL input_rsc_rdy_n_block1_bud : STD_LOGIC;
  SIGNAL output_rsc_vld_n_block1_bud : STD_LOGIC;
  SIGNAL din_rsc_rdy_n_block2_bud : STD_LOGIC;
  SIGNAL dout_rsc_vld_n_block2_bud : STD_LOGIC;

  COMPONENT fir
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      input_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      input_rsc_vld : IN STD_LOGIC;
      input_rsc_rdy : OUT STD_LOGIC;
      coeffs : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      output_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      output_rsc_vld : OUT STD_LOGIC;
      output_rsc_rdy : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL block0_input_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL block0_coeffs : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL block0_output_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);

  SIGNAL block1_input_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL block1_coeffs : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL block1_output_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);

  COMPONENT decimator
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      din_rsc_dat : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      din_rsc_vld : IN STD_LOGIC;
      din_rsc_rdy : OUT STD_LOGIC;
      dout_rsc_dat : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      dout_rsc_vld : OUT STD_LOGIC;
      dout_rsc_rdy : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL block2_din_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL block2_dout_rsc_dat : STD_LOGIC_VECTOR (7 DOWNTO 0);

BEGIN
  block0 : fir
    PORT MAP(
      clk => clk,
      rst => rst,
      input_rsc_dat => block0_input_rsc_dat,
      input_rsc_vld => din_rsc_vld,
      input_rsc_rdy => input_rsc_rdy_n_block0_bud,
      coeffs => block0_coeffs,
      output_rsc_dat => block0_output_rsc_dat,
      output_rsc_vld => output_rsc_vld_n_block0_bud,
      output_rsc_rdy => input_rsc_rdy_n_block1_bud
    );
  block0_input_rsc_dat <= din_rsc_dat;
  block0_coeffs <= coeffs;
  output_rsc_dat_n_block0 <= block0_output_rsc_dat;

  block1 : fir
    PORT MAP(
      clk => clk,
      rst => rst,
      input_rsc_dat => block1_input_rsc_dat,
      input_rsc_vld => output_rsc_vld_n_block0_bud,
      input_rsc_rdy => input_rsc_rdy_n_block1_bud,
      coeffs => block1_coeffs,
      output_rsc_dat => block1_output_rsc_dat,
      output_rsc_vld => output_rsc_vld_n_block1_bud,
      output_rsc_rdy => din_rsc_rdy_n_block2_bud
    );
  block1_input_rsc_dat <= output_rsc_dat_n_block0;
  block1_coeffs <= coeffs;
  output_rsc_dat_n_block1 <= block1_output_rsc_dat;

  block2 : decimator
    PORT MAP(
      clk => clk,
      rst => rst,
      din_rsc_dat => block2_din_rsc_dat,
      din_rsc_vld => output_rsc_vld_n_block1_bud,
      din_rsc_rdy => din_rsc_rdy_n_block2_bud,
      dout_rsc_dat => block2_dout_rsc_dat,
      dout_rsc_vld => dout_rsc_vld_n_block2_bud,
      dout_rsc_rdy => dout_rsc_rdy
    );
  block2_din_rsc_dat <= output_rsc_dat_n_block1;
  dout_rsc_dat_n_block2 <= block2_dout_rsc_dat;

  din_rsc_rdy <= input_rsc_rdy_n_block0_bud;
  dout_rsc_vld <= dout_rsc_vld_n_block2_bud;
  dout_rsc_dat <= dout_rsc_dat_n_block2;
END v2;



